magic
tech sky130A
magscale 1 2
timestamp 1672443751
<< nwell >>
rect 1066 77509 78882 77830
rect 1066 76421 78882 76987
rect 1066 75333 78882 75899
rect 1066 74245 78882 74811
rect 1066 73157 78882 73723
rect 1066 72069 78882 72635
rect 1066 70981 78882 71547
rect 1066 69893 78882 70459
rect 1066 68805 78882 69371
rect 1066 67717 78882 68283
rect 1066 66629 78882 67195
rect 1066 65541 78882 66107
rect 1066 64453 78882 65019
rect 1066 63365 78882 63931
rect 1066 62277 78882 62843
rect 1066 61189 78882 61755
rect 1066 60101 78882 60667
rect 1066 59013 78882 59579
rect 1066 57925 78882 58491
rect 1066 56837 78882 57403
rect 1066 55749 78882 56315
rect 1066 54661 78882 55227
rect 1066 53573 78882 54139
rect 1066 52485 78882 53051
rect 1066 51397 78882 51963
rect 1066 50309 78882 50875
rect 1066 49221 78882 49787
rect 1066 48133 78882 48699
rect 1066 47045 78882 47611
rect 1066 45957 78882 46523
rect 1066 44869 78882 45435
rect 1066 43781 78882 44347
rect 1066 42693 78882 43259
rect 1066 41605 78882 42171
rect 1066 40517 78882 41083
rect 1066 39429 78882 39995
rect 1066 38341 78882 38907
rect 1066 37253 78882 37819
rect 1066 36165 78882 36731
rect 1066 35077 78882 35643
rect 1066 33989 78882 34555
rect 1066 32901 78882 33467
rect 1066 31813 78882 32379
rect 1066 30725 78882 31291
rect 1066 29637 78882 30203
rect 1066 28549 78882 29115
rect 1066 27461 78882 28027
rect 1066 26373 78882 26939
rect 1066 25285 78882 25851
rect 1066 24197 78882 24763
rect 1066 23109 78882 23675
rect 1066 22021 78882 22587
rect 1066 20933 78882 21499
rect 1066 19845 78882 20411
rect 1066 18757 78882 19323
rect 1066 17669 78882 18235
rect 1066 16581 78882 17147
rect 1066 15493 78882 16059
rect 1066 14405 78882 14971
rect 1066 13317 78882 13883
rect 1066 12229 78882 12795
rect 1066 11141 78882 11707
rect 1066 10053 78882 10619
rect 1066 8965 78882 9531
rect 1066 7877 78882 8443
rect 1066 6789 78882 7355
rect 1066 5701 78882 6267
rect 1066 4613 78882 5179
rect 1066 3525 78882 4091
rect 1066 2437 78882 3003
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 1104 1640 78844 77840
<< metal2 >>
rect 39946 79200 40002 80000
rect 1398 0 1454 800
rect 3882 0 3938 800
rect 6366 0 6422 800
rect 8850 0 8906 800
rect 11334 0 11390 800
rect 13818 0 13874 800
rect 16302 0 16358 800
rect 18786 0 18842 800
rect 21270 0 21326 800
rect 23754 0 23810 800
rect 26238 0 26294 800
rect 28722 0 28778 800
rect 31206 0 31262 800
rect 33690 0 33746 800
rect 36174 0 36230 800
rect 38658 0 38714 800
rect 41142 0 41198 800
rect 43626 0 43682 800
rect 46110 0 46166 800
rect 48594 0 48650 800
rect 51078 0 51134 800
rect 53562 0 53618 800
rect 56046 0 56102 800
rect 58530 0 58586 800
rect 61014 0 61070 800
rect 63498 0 63554 800
rect 65982 0 66038 800
rect 68466 0 68522 800
rect 70950 0 71006 800
rect 73434 0 73490 800
rect 75918 0 75974 800
rect 78402 0 78458 800
<< obsm2 >>
rect 1400 79144 39890 79200
rect 40058 79144 78456 79200
rect 1400 856 78456 79144
rect 1510 800 3826 856
rect 3994 800 6310 856
rect 6478 800 8794 856
rect 8962 800 11278 856
rect 11446 800 13762 856
rect 13930 800 16246 856
rect 16414 800 18730 856
rect 18898 800 21214 856
rect 21382 800 23698 856
rect 23866 800 26182 856
rect 26350 800 28666 856
rect 28834 800 31150 856
rect 31318 800 33634 856
rect 33802 800 36118 856
rect 36286 800 38602 856
rect 38770 800 41086 856
rect 41254 800 43570 856
rect 43738 800 46054 856
rect 46222 800 48538 856
rect 48706 800 51022 856
rect 51190 800 53506 856
rect 53674 800 55990 856
rect 56158 800 58474 856
rect 58642 800 60958 856
rect 61126 800 63442 856
rect 63610 800 65926 856
rect 66094 800 68410 856
rect 68578 800 70894 856
rect 71062 800 73378 856
rect 73546 800 75862 856
rect 76030 800 78346 856
<< obsm3 >>
rect 4210 2143 65966 77825
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< labels >>
rlabel metal2 s 41142 0 41198 800 6 a[0]
port 1 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 a[1]
port 2 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 a[2]
port 3 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 a[3]
port 4 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 a[4]
port 5 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 a[5]
port 6 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 a[6]
port 7 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 a[7]
port 8 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 b[0]
port 9 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 b[1]
port 10 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 b[2]
port 11 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 b[3]
port 12 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 b[4]
port 13 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 b[5]
port 14 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 b[6]
port 15 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 b[7]
port 16 nsew signal input
rlabel metal2 s 39946 79200 40002 80000 6 enable
port 17 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 out[0]
port 18 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 out[10]
port 19 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 out[11]
port 20 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 out[12]
port 21 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 out[13]
port 22 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 out[14]
port 23 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 out[15]
port 24 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 out[1]
port 25 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 out[2]
port 26 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 out[3]
port 27 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 out[4]
port 28 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 out[5]
port 29 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 out[6]
port 30 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 out[7]
port 31 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 out[8]
port 32 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 out[9]
port 33 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2811414
string GDS_FILE /home/radhe/shuttle/caravel_user_project/openlane/dadda_multiplier/runs/22_12_31_05_08/results/signoff/dadda_multiplier.magic.gds
string GDS_START 317248
<< end >>

