VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dadda_multiplier
  CLASS BLOCK ;
  FOREIGN dadda_multiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END b[7]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 396.000 200.010 400.000 ;
    END
  END enable
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END out[15]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 387.545 394.410 389.150 ;
        RECT 5.330 382.105 394.410 384.935 ;
        RECT 5.330 376.665 394.410 379.495 ;
        RECT 5.330 371.225 394.410 374.055 ;
        RECT 5.330 365.785 394.410 368.615 ;
        RECT 5.330 360.345 394.410 363.175 ;
        RECT 5.330 354.905 394.410 357.735 ;
        RECT 5.330 349.465 394.410 352.295 ;
        RECT 5.330 344.025 394.410 346.855 ;
        RECT 5.330 338.585 394.410 341.415 ;
        RECT 5.330 333.145 394.410 335.975 ;
        RECT 5.330 327.705 394.410 330.535 ;
        RECT 5.330 322.265 394.410 325.095 ;
        RECT 5.330 316.825 394.410 319.655 ;
        RECT 5.330 311.385 394.410 314.215 ;
        RECT 5.330 305.945 394.410 308.775 ;
        RECT 5.330 300.505 394.410 303.335 ;
        RECT 5.330 295.065 394.410 297.895 ;
        RECT 5.330 289.625 394.410 292.455 ;
        RECT 5.330 284.185 394.410 287.015 ;
        RECT 5.330 278.745 394.410 281.575 ;
        RECT 5.330 273.305 394.410 276.135 ;
        RECT 5.330 267.865 394.410 270.695 ;
        RECT 5.330 262.425 394.410 265.255 ;
        RECT 5.330 256.985 394.410 259.815 ;
        RECT 5.330 251.545 394.410 254.375 ;
        RECT 5.330 246.105 394.410 248.935 ;
        RECT 5.330 240.665 394.410 243.495 ;
        RECT 5.330 235.225 394.410 238.055 ;
        RECT 5.330 229.785 394.410 232.615 ;
        RECT 5.330 224.345 394.410 227.175 ;
        RECT 5.330 218.905 394.410 221.735 ;
        RECT 5.330 213.465 394.410 216.295 ;
        RECT 5.330 208.025 394.410 210.855 ;
        RECT 5.330 202.585 394.410 205.415 ;
        RECT 5.330 197.145 394.410 199.975 ;
        RECT 5.330 191.705 394.410 194.535 ;
        RECT 5.330 186.265 394.410 189.095 ;
        RECT 5.330 180.825 394.410 183.655 ;
        RECT 5.330 175.385 394.410 178.215 ;
        RECT 5.330 169.945 394.410 172.775 ;
        RECT 5.330 164.505 394.410 167.335 ;
        RECT 5.330 159.065 394.410 161.895 ;
        RECT 5.330 153.625 394.410 156.455 ;
        RECT 5.330 148.185 394.410 151.015 ;
        RECT 5.330 142.745 394.410 145.575 ;
        RECT 5.330 137.305 394.410 140.135 ;
        RECT 5.330 131.865 394.410 134.695 ;
        RECT 5.330 126.425 394.410 129.255 ;
        RECT 5.330 120.985 394.410 123.815 ;
        RECT 5.330 115.545 394.410 118.375 ;
        RECT 5.330 110.105 394.410 112.935 ;
        RECT 5.330 104.665 394.410 107.495 ;
        RECT 5.330 99.225 394.410 102.055 ;
        RECT 5.330 93.785 394.410 96.615 ;
        RECT 5.330 88.345 394.410 91.175 ;
        RECT 5.330 82.905 394.410 85.735 ;
        RECT 5.330 77.465 394.410 80.295 ;
        RECT 5.330 72.025 394.410 74.855 ;
        RECT 5.330 66.585 394.410 69.415 ;
        RECT 5.330 61.145 394.410 63.975 ;
        RECT 5.330 55.705 394.410 58.535 ;
        RECT 5.330 50.265 394.410 53.095 ;
        RECT 5.330 44.825 394.410 47.655 ;
        RECT 5.330 39.385 394.410 42.215 ;
        RECT 5.330 33.945 394.410 36.775 ;
        RECT 5.330 28.505 394.410 31.335 ;
        RECT 5.330 23.065 394.410 25.895 ;
        RECT 5.330 17.625 394.410 20.455 ;
        RECT 5.330 12.185 394.410 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 5.520 8.200 394.220 389.200 ;
      LAYER met2 ;
        RECT 7.000 395.720 199.450 396.000 ;
        RECT 200.290 395.720 392.280 396.000 ;
        RECT 7.000 4.280 392.280 395.720 ;
        RECT 7.550 4.000 19.130 4.280 ;
        RECT 19.970 4.000 31.550 4.280 ;
        RECT 32.390 4.000 43.970 4.280 ;
        RECT 44.810 4.000 56.390 4.280 ;
        RECT 57.230 4.000 68.810 4.280 ;
        RECT 69.650 4.000 81.230 4.280 ;
        RECT 82.070 4.000 93.650 4.280 ;
        RECT 94.490 4.000 106.070 4.280 ;
        RECT 106.910 4.000 118.490 4.280 ;
        RECT 119.330 4.000 130.910 4.280 ;
        RECT 131.750 4.000 143.330 4.280 ;
        RECT 144.170 4.000 155.750 4.280 ;
        RECT 156.590 4.000 168.170 4.280 ;
        RECT 169.010 4.000 180.590 4.280 ;
        RECT 181.430 4.000 193.010 4.280 ;
        RECT 193.850 4.000 205.430 4.280 ;
        RECT 206.270 4.000 217.850 4.280 ;
        RECT 218.690 4.000 230.270 4.280 ;
        RECT 231.110 4.000 242.690 4.280 ;
        RECT 243.530 4.000 255.110 4.280 ;
        RECT 255.950 4.000 267.530 4.280 ;
        RECT 268.370 4.000 279.950 4.280 ;
        RECT 280.790 4.000 292.370 4.280 ;
        RECT 293.210 4.000 304.790 4.280 ;
        RECT 305.630 4.000 317.210 4.280 ;
        RECT 318.050 4.000 329.630 4.280 ;
        RECT 330.470 4.000 342.050 4.280 ;
        RECT 342.890 4.000 354.470 4.280 ;
        RECT 355.310 4.000 366.890 4.280 ;
        RECT 367.730 4.000 379.310 4.280 ;
        RECT 380.150 4.000 391.730 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 329.830 389.125 ;
  END
END dadda_multiplier
END LIBRARY

